*
vin	Vin	0	AC	1V
*
C6	Vin	1	0.1u
R4	1	2	10K
D1	2	0	1N4148
D2	0	2	1N4148
R6	2	3	6.8k
C8	3	4	0.022u
R5	4	0	1k
C9	3	5	0.22u
P1	4	5	5	100k
C7	2	6	0.022u
P2	5	vout	5	22k
*
*	V-	V+	out
Z2a	4	2	vout

.MODEL 1N4148 D (IS=4.352e-9 N=1.906 BV=110 IBV=0.0001 RS=0.6458 CJO=7.048e-13 VJ=0.869 M=0.03 FC=0.5 TT=3.48e-9)
